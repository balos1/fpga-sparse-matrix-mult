/*
    Test bench for communication module.

    author(s): Cody Balos <cjbalos@gmail.com>
*/

module test_comm_unit();




endmodule
